StudentSenseHatV06
R4 3 7 3.9k
R7 1 5 4.7k
R1 4 8 1k
R9 4 8 1k
R5 3 2 3.9k
R6 1 6 4.7k

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
